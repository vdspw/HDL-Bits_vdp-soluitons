//Problem : Build a circuit with no inputs and one output that outputs a constant 0


module top_module(
    output zero
);
assign zero = 1'b0;
// Output data type is used and variable zero is declared.
// using assign statement the output is driven.
endmodule
